package MAL is 
 	 component place_b 
 	 	 port(ck, ra0_int, ra1_init, activer, desactiver : in std_logic ;
 	 	 	 marque : out std_logic) ;
 	end component ; 
end MAL ;

